`timescale 1ns / 1ps
`include "riscv_define.v"

module MemorySystem_tb;

    // === 1. �źŶ��� ===
    reg clk;
    reg rst_n;
    reg flush;

    // LSU (D-Cache) �����ź�
    reg lsu_valid_in;
    reg [31:0] lsu_addr;
    reg [31:0] lsu_wdata;
    reg [`MEM_OP_WIDTH-1:0] lsu_op;
    reg lsu_is_load;
    reg lsu_unsigned;
    
    // LSU ����۲�
    wire lsu_busy;
    wire lsu_wb_valid;
    wire [31:0] lsu_wb_value;

    // I-Cache �����ź�
    reg [31:0] if_pc;
    reg if_req;
    
    // I-Cache ����۲�
    wire [127:0] if_inst_line;
    wire if_hit;
    wire if_stall;

    // �ڲ������ź� (Arbiter <-> Memory)
    wire arb_mem_req, arb_mem_we, arb_mem_ready;
    wire [31:0] arb_mem_addr;
    wire [127:0] arb_mem_wdata, arb_mem_rdata;

    // �����ź� (Components <-> Arbiter)
    wire i_req, i_we, i_ready;
    wire [31:0] i_addr;
    wire [127:0] i_wdata, i_rdata;
    
    wire d_req, d_we, d_ready;
    wire [31:0] d_addr;
    wire [127:0] d_wdata, d_rdata;

    // === 2. ģ��ʵ���� ===

    // 2.1 ������ģ�LSU (�� TLB + D-Cache)
    LSU u_lsu (
        .clk(clk), .rst_n(rst_n), .flush(flush),
        .valid_in(lsu_valid_in),
        .addr(lsu_addr),
        .wdata(lsu_wdata),
        .mem_op(lsu_op),
        .mem_is_load(lsu_is_load),
        .mem_unsigned(lsu_unsigned),
        .rob_idx_in(0), .rd_tag_in(1), .rd_is_fp_in(0), // �򵥵� dummy �ź�
        .busy(lsu_busy),
        .wb_valid(lsu_wb_valid),
        .wb_value(lsu_wb_value),
        // ���ӵ� Arbiter �� D �˿�
        .mem_req(d_req), .mem_we(d_we), .mem_addr(d_addr),
        .mem_wdata(d_wdata), .mem_rdata(d_rdata), .mem_ready(d_ready)
    );

    // 2.2 ������ģ�ICache
    ICache u_icache (
        .clk(clk), .rst_n(rst_n),
        .paddr(if_pc),
        .req(if_req),
        .rdata_line(if_inst_line),
        .valid_out(if_hit),
        .stall_cpu(if_stall),
        // ���ӵ� Arbiter �� I �˿�
        .mem_req(i_req), .mem_we(i_we), .mem_addr(i_addr),
        .mem_wdata(i_wdata), .mem_rdata(i_rdata), .mem_ready(i_ready)
    );

    // 2.3 �ٲ���
    MemArbiter u_arbiter (
        .clk(clk), .rst_n(rst_n),
        .i_req(i_req), .i_we(i_we), .i_addr(i_addr), .i_wdata(i_wdata), .i_rdata(i_rdata), .i_ready(i_ready),
        .d_req(d_req), .d_we(d_we), .d_addr(d_addr), .d_wdata(d_wdata), .d_rdata(d_rdata), .d_ready(d_ready),
        .mem_req(arb_mem_req), .mem_we(arb_mem_we), .mem_addr(arb_mem_addr), .mem_wdata(arb_mem_wdata), .mem_rdata(arb_mem_rdata), .mem_ready(arb_mem_ready)
    );

    // 2.4 ����ģ��
    MainMemory u_mem (
        .clk(clk), .rst_n(rst_n),
        .mem_req(arb_mem_req), .mem_we(arb_mem_we), .mem_addr(arb_mem_addr), .mem_wdata(arb_mem_wdata),
        .mem_rdata(arb_mem_rdata), .mem_ready(arb_mem_ready)
    );

    // === 3. ʱ������ ===
    always #5 clk = ~clk; // 100MHz

    // === 4. �������� (Helper Tasks) ===
    
    // ���񣺸�λ
    task reset_system;
    begin
        $display("\n[TEST] System Reset...");
        clk = 0; rst_n = 0; flush = 0;
        lsu_valid_in = 0; if_req = 0;
        #20 rst_n = 1;
        #10;
    end
    endtask

    // ����LSU Store
    task lsu_store(input [31:0] addr, input [31:0] data);
    begin
        $display("[LSU] STORE Request: Addr=0x%h, Data=0x%h", addr, data);
        @(posedge clk);
        lsu_valid_in = 1;
        lsu_addr = addr;
        lsu_wdata = data;
        lsu_op = `MEM_OP_SW;
        lsu_is_load = 0;
        
        // �ȴ� Busy
        @(posedge clk);
        lsu_valid_in = 0;
        
        // �ȴ���� (wb_valid ���� Store Ҳ������Ϊ��ɱ�־�����߿� busy ���)
        wait(lsu_wb_valid);
        $display("[LSU] STORE Completed.");
        @(posedge clk);
    end
    endtask

    // ����LSU Load
    task lsu_load(input [31:0] addr, input [31:0] expected_data);
    begin
        $display("[LSU] LOAD Request:  Addr=0x%h", addr);
        @(posedge clk);
        lsu_valid_in = 1;
        lsu_addr = addr;
        lsu_op = `MEM_OP_LW;
        lsu_is_load = 1;
        
        @(posedge clk);
        lsu_valid_in = 0;
        
        wait(lsu_wb_valid);
        if (lsu_wb_value === expected_data) 
            $display("[PASS] LSU Load Hit/Miss Success! Got 0x%h", lsu_wb_value);
        else 
            $display("[FAIL] LSU Load Error! Expected 0x%h, Got 0x%h", expected_data, lsu_wb_value);
        @(posedge clk);
    end
    endtask

    // ����ICache Fetch
    task icache_fetch(input [31:0] addr);
    begin
        $display("[IF]  FETCH Request: Addr=0x%h", addr);
        @(posedge clk);
        if_pc = addr;
        if_req = 1;
        
        // �ȴ� valid_out (Hit)
        // ע�⣺����� Miss��valid_out �����������ں���
        wait(if_hit); 
        $display("[PASS] ICache Valid! Data Line: 0x%h", if_inst_line);
        if_req = 0; // ֹͣ����
        @(posedge clk);
    end
    endtask

    // === 5. ���������� ===
    initial begin
        // ��ʼ���������� (�� MainMemory.v ��ͨ������ initial block�������������)
        // �����ַ 0x00 ���������� 0xDEAD_BEEF... (��� MainMemory.v д��)

        reset_system();

        // --- Test 1: I-Cache Cold Miss (��һ�ζ�) ---
        $display("\n--- Test 1: I-Cache Cold Miss ---");
        // �����ַ 0 ��Ӧ Set 0
        icache_fetch(32'h0000_0000); 

        // --- Test 2: I-Cache Hit (�ڶ��ζ�ͬһ��ַ) ---
        $display("\n--- Test 2: I-Cache Hit ---");
        // Ӧ���� 1 �������ڷ��ؽ��������Ҫ arbiter ����
        icache_fetch(32'h0000_0004); // ͬһ�� Cache Line��Ӧ��ֱ�� Hit

        // --- Test 3: LSU Store (д�� D-Cache) ---
        $display("\n--- Test 3: LSU Store ---");
        // ����ַ 0x100 д�� 0x12345678
        lsu_store(32'h0000_0100, 32'h1234_5678);

        // --- Test 4: LSU Load (��ȡ�ղ�д�������) ---
        $display("\n--- Test 4: LSU Load (Read after Write) ---");
        // �ӵ�ַ 0x100 ����Ӧ������ D-Cache ������ 0x12345678
        lsu_load(32'h0000_0100, 32'h1234_5678);

        // --- Test 5: Conflict Test (ICache Miss + LSU Miss) ---
        $display("\n--- Test 5: Conflict Test (Arbiter) ---");
        $display("[TEST] Asserting both requests simultaneously...");
        
        @(posedge clk);
        // ����һ���µ� Miss
        if_pc = 32'h0000_0200; if_req = 1; // I-Cache ����
        
        lsu_valid_in = 1; lsu_addr = 32'h0000_0300; lsu_op = `MEM_OP_LW; lsu_is_load = 1; // LSU ����
        
        @(posedge clk);
        lsu_valid_in = 0; // LSU �������ź�
        // if_req ���ָߵ�ƽֱ�� hit
        
        $display("[TEST] Waiting for completion...");
        
        // ����������ɣ�˳��ȡ���� Arbiter (����� D ����)
        fork
            begin
                wait(lsu_wb_valid);
                $display("[INFO] LSU Finished first (Expected behavior).");
            end
            begin
                wait(if_hit);
                $display("[INFO] ICache Finished.");
            end
        join

        $display("\n[SUCCESS] All Tests Passed!");
        $finish;
    end

    // ��� Arbiter ״̬ (������)
    always @(posedge clk) begin
        if (arb_mem_req && arb_mem_ready)
            $display("    [MEM] Transaction Addr=0x%h Data=0x%h", arb_mem_addr, arb_mem_rdata);
    end

endmodule