// ram.v
module ram #(
    parameter ADDR_WIDTH = 12,   // RAM ��� = 2^ADDR_WIDTH
    parameter DATA_WIDTH = 32
)(
    input  wire                   clk,

    // д�˿ڣ�����д�� dirty �У�
    input  wire                   we,
    input  wire [ADDR_WIDTH-1:0]  waddr,
    input  wire [DATA_WIDTH-1:0]  din,

    // ���˿ڣ����ڶ� miss ʱ���ڴ�ȡ���ݣ�
    input  wire [ADDR_WIDTH-1:0]  raddr,
    output wire [DATA_WIDTH-1:0]  dout
);

    localparam DEPTH = 1 << ADDR_WIDTH;

    reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];

    // д��ͬ��
    always @(posedge clk) begin
        if (we)
            mem[waddr] <= din;
    end

    // ������ϣ���ѧ�Ѻã����ӳ٣�
    assign dout = mem[raddr];

endmodule
