// cache_and_ram.v
module cache_and_ram #(
    parameter ADDR_WIDTH  = 12,       // ���� cache �ĵ�ַλ��
    parameter INDEX_WIDTH = 6,        // ���λ�� -> ���� = 2^INDEX_WIDTH
    parameter DATA_WIDTH  = 32
)(
    input  wire                   clk,
    input  wire                   rst,

    input  wire                   mode,        // 1 = write, 0 = read
    input  wire [31:0]            address,     // CPU �ӽǵ�ַ��ֻ�õ� ADDR_WIDTH λ��
    input  wire [DATA_WIDTH-1:0]  data_in,     // CPU д����

    output reg  [DATA_WIDTH-1:0]  out,         // CPU ������
    output reg                    out_valid    // �������Ƿ���Ч
);

    // ------------------------------
    // ��ַ��֣��� INDEX_WIDTH λ�� index���� TAG_WIDTH λ�� tag
    // ------------------------------
    localparam TAG_WIDTH = ADDR_WIDTH - INDEX_WIDTH;
    localparam LINE_NUM  = 1 << INDEX_WIDTH;

    wire [ADDR_WIDTH-1:0]  addr_in   = address[ADDR_WIDTH-1:0];
    wire [INDEX_WIDTH-1:0] index     = addr_in[INDEX_WIDTH-1:0];
    wire [TAG_WIDTH-1:0]   tag       = addr_in[ADDR_WIDTH-1:INDEX_WIDTH];

    // ���� RAM ����ȡ�¿飩
    wire [ADDR_WIDTH-1:0]  ram_raddr = addr_in;

    // ------------------------------
    // �滻���ԣ�ÿ��һ�� bit��0 ��ʾѡ way0��1 ��ʾѡ way1
    // ����ת���൱��ÿ��� random / round-robin
    // ------------------------------
    reg repl_bit [0:LINE_NUM-1];

    integer k;
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            for (k = 0; k < LINE_NUM; k = k + 1)
                repl_bit[k] <= 1'b0;
        end else begin
            // �� miss ʱ�ŷ�ת repl_bit[index]�������߼���ʵ��
        end
    end

    // ��ϳ���ǰ����滻��ѡ way
    wire [0:0] evict_way = repl_bit[index];

    // ------------------------------
    // Cache 2-way ʵ��
    // ------------------------------
    wire        cache_hit;
    wire [0:0]  cache_hit_way;
    wire [DATA_WIDTH-1:0] cache_dout;

    reg         cache_we;
    reg  [0:0]  cache_way_sel;
    reg  [DATA_WIDTH-1:0] cache_din;
    reg         cache_valid_in;
    reg         cache_dirty_in;

    wire        sel_valid;
    wire        sel_dirty;
    wire [TAG_WIDTH-1:0]   sel_tag;
    wire [DATA_WIDTH-1:0]  sel_data;

    cache_2way #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .TAG_WIDTH  (TAG_WIDTH),
        .DATA_WIDTH (DATA_WIDTH),
        .WAYS       (2)
    ) u_cache (
        .clk       (clk),
        .rst       (rst),
        .index     (index),
        .tag_in    (tag),
        .we        (cache_we),
        .way_sel   (cache_way_sel),
        .din       (cache_din),
        .valid_in  (cache_valid_in),
        .dirty_in  (cache_dirty_in),
        .hit       (cache_hit),
        .hit_way   (cache_hit_way),
        .dout      (cache_dout),
        .sel_valid (sel_valid),
        .sel_dirty (sel_dirty),
        .sel_tag   (sel_tag),
        .sel_data  (sel_data)
    );

    // ------------------------------
    // RAM ʵ����һдһ��
    // д�˿����� write-back�����˿����� miss refill
    // ------------------------------
    reg                  ram_we;
    reg  [ADDR_WIDTH-1:0] ram_waddr;
    reg  [DATA_WIDTH-1:0] ram_din;
    wire [DATA_WIDTH-1:0] ram_dout;

    ram #(
        .ADDR_WIDTH(ADDR_WIDTH),
        .DATA_WIDTH(DATA_WIDTH)
    ) u_ram (
        .clk   (clk),
        .we    (ram_we),
        .waddr (ram_waddr),
        .din   (ram_din),
        .raddr (ram_raddr),
        .dout  (ram_dout)
    );

    // ------------------------------
    // �������߼�
    // д���ԣ�д�� + д����
    // �滻���ԣ�ÿ���ֻ� evict_way
    // ------------------------------
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            out       <= {DATA_WIDTH{1'b0}};
            out_valid <= 1'b0;

            cache_we       <= 1'b0;
            cache_way_sel  <= 1'b0;
            cache_din      <= {DATA_WIDTH{1'b0}};
            cache_valid_in <= 1'b0;
            cache_dirty_in <= 1'b0;

            ram_we    <= 1'b0;
            ram_waddr <= {ADDR_WIDTH{1'b0}};
            ram_din   <= {DATA_WIDTH{1'b0}};
        end else begin
            // Ĭ�ϲ�д cache / ram
            cache_we       <= 1'b0;
            cache_valid_in <= 1'b0;
            cache_dirty_in <= 1'b0;
            ram_we         <= 1'b0;
            out_valid      <= 1'b0;

            // ѡ�ĸ� way��д����ʱѡ�� hit_way������ѡ�� evict_way
            cache_way_sel <= (cache_hit && mode) ? cache_hit_way : evict_way;

            if (mode) begin
                //--------------------------------------
                // д������write-back + write-allocate
                //--------------------------------------
                if (cache_hit) begin
                    // д���У�ֻд cache����Ӧ�� dirty=1��������д RAM
                    cache_we       <= 1'b1;
                    cache_din      <= data_in;
                    cache_valid_in <= 1'b1;
                    cache_dirty_in <= 1'b1;    // д�ز��ԣ����Ϊ dirty

                    // ��д RAM��д�أ�
                    ram_we         <= 1'b0;
                end else begin
                    // д miss��д���䣨write-allocate��
                    // 1) ���滻���� valid �� dirty����Ҫд��
                    if (sel_valid && sel_dirty) begin
                        ram_we    <= 1'b1;
                        ram_waddr <= {sel_tag, index};  // �ñ��滻�е� tag + index ��ԭ��ַ
                        ram_din   <= sel_data;          // д�ؾ�����
                    end

                    // 2) �� cache �з������У�ֱ��д�� data_in������� dirty
                    cache_we       <= 1'b1;
                    cache_din      <= data_in;
                    cache_valid_in <= 1'b1;
                    cache_dirty_in <= 1'b1;  // д���� dirty

                    // 3) �����滻λ�������ֻ��´��滻�� way
                    repl_bit[index] <= ~repl_bit[index];

                    // д����һ�㲻�� CPU ��������
                    out_valid <= 1'b0;
                end

            end else begin
                //--------------------------------------
                // ������
                //--------------------------------------
                if (cache_hit) begin
                    // �����У�ֱ�Ӵ� cache ȡ����
                    out       <= cache_dout;
                    out_valid <= 1'b1;

                    // ����Ҫд RAM / cache
                end else begin
                    // �� miss����Ҫ�� RAM ȡ���ݣ�������д�ر��滻 dirty ��

                    // 1) ������滻�� dirty����д��
                    if (sel_valid && sel_dirty) begin
                        ram_we    <= 1'b1;
                        ram_waddr <= {sel_tag, index};
                        ram_din   <= sel_data;
                    end

                    // 2) �� RAM �������ݣ�ram_dout �Ѿ��� raddr ��Ӧ��ֵ��
                    //    д�� cache��valid=1, dirty=0����Ϊ�Ǵ��ڴ�ն����ĸɾ����ݣ�
                    cache_we       <= 1'b1;
                    cache_din      <= ram_dout;
                    cache_valid_in <= 1'b1;
                    cache_dirty_in <= 1'b0;  // fresh from memory

                    // 3) ���ظ� CPU
                    out       <= ram_dout;
                    out_valid <= 1'b1;

                    // 4) ���¸�����滻��Ϣ
                    repl_bit[index] <= ~repl_bit[index];
                end
            end
        end
    end

endmodule
