// simple_tlb.v
module tlb #(
    parameter ENTRY_NUM = 16,        // TLB ��������
    parameter VPN_WIDTH = 20,        // ����ҳ��λ��Sv32: 32-12=20��
    parameter PPN_WIDTH = 20         // ����ҳ��λ��
)(
    input  wire                  clk,
    input  wire                  rst,

    // ========= ���ӿڣ��� MEM / cache �ã� =========
    input  wire [31:0]           lookup_vaddr,   // �����ַ
    output wire [31:0]           lookup_paddr,   // �����ַ������ʱ��Ч��
    output wire                  lookup_hit,     // �Ƿ�����
    output wire                  lookup_pagefault, // ҳ�쳣�����������ӿڣ�һ�� 0��

    // ========= д��ӿڣ��Ժ� OS ͨ����Ȩָ�����ã� =========
    input  wire                  wr_en,          // д��һ�� TLB ����
    input  wire [31:0]           wr_vaddr,       // ��Ӧ�����ַ��ֻ�� VPN ���֣�
    input  wire [31:0]           wr_paddr,       // ��Ӧ�����ַ��ֻ�� PPN ���֣�
    input  wire [2:0]            wr_perm,        // Ȩ�ޱ�־��R/W/X�����ڲ�ϸ�ã��ȴ��ţ�

    // ========= ˢ�½ӿڣ�sfence.vma ֮�ࣩ =========
    input  wire                  flush           // �� 1 ʱ������� TLB ����
);

    // ---- TLB ����洢 ----
    reg                  valid   [0:ENTRY_NUM-1];
    reg [VPN_WIDTH-1:0]  vpn     [0:ENTRY_NUM-1];
    reg [PPN_WIDTH-1:0]  ppn     [0:ENTRY_NUM-1];
    reg [2:0]            perm    [0:ENTRY_NUM-1]; // �ȴ�������������Ȩ��У����

    // �� round-robin �滻ָ��
    reg [$clog2(ENTRY_NUM)-1:0] rr_ptr;

    integer i;

    // ---- ����߼���ȫ�������� ----
    wire [VPN_WIDTH-1:0] curr_vpn   = lookup_vaddr[31:32-VPN_WIDTH];
    wire [11:0]          page_off   = lookup_vaddr[11:0];

    reg                  hit_r;
    reg [PPN_WIDTH-1:0]  hit_ppn;

    always @(*) begin
        hit_r   = 1'b0;
        hit_ppn = {PPN_WIDTH{1'b0}};
        for (i = 0; i < ENTRY_NUM; i = i + 1) begin
            if (valid[i] && vpn[i] == curr_vpn) begin
                hit_r   = 1'b1;
                hit_ppn = ppn[i];
            end
        end
    end

    assign lookup_hit        = hit_r;
    assign lookup_paddr      = {hit_ppn, page_off};
    assign lookup_pagefault  = 1'b0;   // �����Ȳ���Ȩ����ҳ��У�飬ͳһ�� 0

    // ---- д�� / �滻�߼� ----
    reg [$clog2(ENTRY_NUM)-1:0] free_idx;
    reg                         has_free;

    // ����û�� invalid �Ŀ�λ����ϣ�
    always @(*) begin
        has_free = 1'b0;
        free_idx = {($clog2(ENTRY_NUM)){1'b0}};
        for (i = 0; i < ENTRY_NUM; i = i + 1) begin
            if (!valid[i]) begin
                has_free = 1'b1;
                free_idx = i[$clog2(ENTRY_NUM)-1:0];
            end
        end
    end

    // ʱ�򲿷֣�reset / flush / wr_en
    integer j;
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            rr_ptr <= {($clog2(ENTRY_NUM)){1'b0}};
            for (j = 0; j < ENTRY_NUM; j = j + 1) begin
                valid[j] <= 1'b0;
                vpn[j]   <= {VPN_WIDTH{1'b0}};
                ppn[j]   <= {PPN_WIDTH{1'b0}};
                perm[j]  <= 3'b000;
            end
        end else begin
            if (flush) begin
                for (j = 0; j < ENTRY_NUM; j = j + 1) begin
                    valid[j] <= 1'b0;
                end
            end else if (wr_en) begin
                // �п�λ��д��λ�������� rr_ptr �滻
                if (has_free) begin
                    valid[free_idx] <= 1'b1;
                    vpn[free_idx]   <= wr_vaddr[31:32-VPN_WIDTH];
                    ppn[free_idx]   <= wr_paddr[31:32-PPN_WIDTH];
                    perm[free_idx]  <= wr_perm;
                end else begin
                    valid[rr_ptr] <= 1'b1;
                    vpn[rr_ptr]   <= wr_vaddr[31:32-VPN_WIDTH];
                    ppn[rr_ptr]   <= wr_paddr[31:32-PPN_WIDTH];
                    perm[rr_ptr]  <= wr_perm;
                    rr_ptr        <= rr_ptr + 1'b1;
                end
            end
        end
    end

endmodule
